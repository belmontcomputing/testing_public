module test_pub;
endmodule
